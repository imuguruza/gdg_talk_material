module top(
            input i_clk,
            input i_en,
            input i_reset,
            output o_tx,
            output o_led);

always @(posedge clk) begin

endmodule
