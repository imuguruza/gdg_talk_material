`define clk	12000000
