//
`define alhambra_clk	12000000
`define ulx3s_clk	12000000
